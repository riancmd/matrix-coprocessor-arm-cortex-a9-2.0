`timescale 1ns / 1ps

module testMultM();
    reg rst;
    reg signed [199:0] lin, col;  // 200 bits => matrizes 5x5
    wire signed [199:0] n_out;    // 200 bits => matriz 5x5
    wire ovf;
    
    // Instância do módulo de multiplicação

    mult_M uut(
        .lin(lin),
        .col(col),
        .rst(rst),
        .n_out(n_out),
        .ovf(ovf)
    );
    
    
    // Gera sinal de reset
    initial begin
        $display("Inicia reset");
        rst = 1'b1;
        #10 rst = 1'b0;
    end
    
    // Testa os estímulos
    initial begin
        $display("Testa valores");
        $monitor("tempo=%3d, rst=%b, lin=%200b, col=%200b, n_out=%200b, ovf=%b", 
                 $time, rst, lin, col, n_out, ovf);
            
        #15; // Espera reset terminar
            
        // CASO 1: Valores pequenos positivos (sem overflow)
        // lin = [1, 2, 3, 4, 2, 1, 2, 1, 2, 3, 1, 2, 1, 1, 2, 2, 2, 1, 3, 2, 2, 1, 1, 2, 2]
        lin = 200'b00000001_00000010_00000011_00000100_00000010_00000001_00000010_00000001_00000010_00000011_00000001_00000010_00000001_00000001_00000010_00000010_00000010_00000001_00000011_00000010_00000010_00000001_00000001_00000010_00000010;
        // col = [ 2, 1, 2, 3, 2, 1, 2, 3, 1, 2, 1, 2, 0, 3, 3, 2, 2, 1, 1, 3, 2, 1, 1, 2, 0] 
        col = 200'b00000010_00000001_00000001_00000010_00000010_00000001_00000010_00000010_00000010_00000001_00000010_00000001_00000001_00000010_00000001_00000011_00000011_00000000_00000001_00000011_00000010_00000010_00000001_00000010_00000000;
        // n_out esperado: [19, 21, 14, 22, 27, 15, 14, 13, 16, 15, 11, 11, 11, 13, 12, 41, 71, 61, 51, 82, 05, 14, 12, 11, 16, 15]
        // Resultado esperado: 200'b00010011_00010101_00001110_00010110_00011011_00001111_00001110_00001101_00010000_00001111_00001011_00001011_00001011_00001101_00001100_00101001_01000111_00111101_00110011_01010010_00000101_00001110_00001100_00001011_00010000;
        
    end
endmodule