module buffer_2x2_HPStoFGPA(
	input [199:0] matrix1_in, matrix2_in, //Matrizes vindo sem organização
	output [199:0] matrix1_out, matrix2_out //Matrizes organizadas com base no tamanho
);
	
	//Organizando a matriz 1
	assign matrix1_out[199:184] = matrix1_in[199:184];
	assign matrix1_out[159:144] = matrix1_in[183:168];
	
	assign matrix1_out[183:160] = 0;
	assign matrix1_out[143:0] = 0;

	
	//Organizando a matriz 2
	assign matrix2_out[199:184] = matrix2_in[199:184];
	assign matrix2_out[159:144] = matrix2_in[183:168];
	
	assign matrix2_out[183:160] = 0;
	assign matrix2_out[143:0] = 0;
	
endmodule